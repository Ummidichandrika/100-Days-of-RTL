//interface
interface fs_if;
logic a;
logic b;
logic bin;
logic diff;
logic bout;
endinterface
