//transaction.sv
class transaction;
randc bit a;
randc bit b; 

bit sum;
bit cout;
endclass
