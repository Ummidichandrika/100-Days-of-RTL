//interface
interface ha_if;
  
logic a;
logic b;
logic sum;
logic cout;
  
endinterface
