class transaction;

  rand bit[3:0] d;
  rand bit  [1:0]    sel;
  bit    y;

  

endclass
