//transaction.sv
class transaction;
randc bit a;
randc bit b;
randc bit bin; 
bit diff;
bit bout;
endclass
