interface mux_if();
  logic [3:0] d;
  logic [1:0] sel;
  logic y;
  
endinterface 
  
