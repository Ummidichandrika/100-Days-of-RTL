//interface
interface dec_if;
  logic [2:0] d;
  logic [7:0] o;

endinterface
