//transaction.sv
class transaction;
  randc bit [2:0] d;
  bit[7:0] o ;

endclass
